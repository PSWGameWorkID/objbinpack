/* SPDX-License-Identifier: GPL-3.0 */
/**
 * maker_c.v
 * 
 * PURPOSE
 *  C code generator and gcc/clang compiler feeder for objbinpack
 * 
 * COPYRIGHT
 *  (C) 2025 Syahriel "EmiyaSyahriel" Ibnu Irfansyah
 */

module main
import os

struct MakerC
{
pub mut:
	cc string
	state States
}

fn (mut this MakerC) process(states States) 
{
	this.cc = os.getenv_opt("CC") or { "gcc" }
	this.cc = os.find_abs_path_of_executable(this.cc) or { os.abs_path(this.cc) }
	mut process := os.new_process(this.cc)
	oflags := parse_oflags(states.cflags)
	mut args := ["-o", states.out_path, "-x", "c", "-c", "-"]
	args << oflags.data
	
	process.set_args(args)
	process.set_redirect_stdio()
	println("MakeC : starting ${this.cc}")
	process.run()
	println("MakeC : ${this.cc} startup success ( PID ${process.pid} ), C writing source header...")
	
	process.stdin_write("/** Generated by objbinpack - no one gonna read it this though since this is directly pushed to compiled via stdin */\r")
	process.stdin_write("#include <stdint.h>\r\n")
	process.stdin_write("#include <stddef.h>\r\n")
	for input in states.inputs {
		println("MakeC : writing \"${input.file_path}\" as \"${input.variable_name}\"")
		varname := input.variable_name 
		fsize := os.file_size(input.file_path)
		process.stdin_write("const uint8_t ${varname}_data[] = {\n\t");
		file := os.open(input.file_path)  or { panic(err) }
		mut bytes_read := 0;
		mut buffer := []u8{len:64}
		for !file.eof() {
			buf_read := file.read(mut buffer) or { panic(err) }
			for i in 0 .. buf_read {
				a_byte := buffer[i]
				process.stdin_write("0x${a_byte.hex()}")
				if bytes_read < fsize - 1 {
					process.stdin_write(",")
				}
				bytes_read++
			}
		}
		
		process.stdin_write("\n};\n")
		process.stdin_write("const size_t ${varname}_length = ${fsize};\n")
	}

	println("MakeC : finishing up")
	os.fd_close(process.stdio_fd[0])
	s_stdout := process.stdout_slurp()
	s_stderr := process.stderr_slurp()
	println("MakeC : waiting for ${this.cc} to exit...")
	process.wait()
	println("${this.cc} STDOUT: ")
	println(s_stdout)
	println("${this.cc} STDERR: ")
	println(s_stderr)
	println("MakeC : ${this.cc} exited with code ${process.code} (${process.err}), cleaning up...")
	process.close()
}