/* SPDX-License-Identifier: GPL-3.0 */
/**
 * maker_cpp.v
 * 
 * PURPOSE
 *  C++ code generator and g++/clang++ compiler feeder for objbinpack
 * 
 * COPYRIGHT
 *  (C) 2025 Syahriel "EmiyaSyahriel" Ibnu Irfansyah
 */

module main
import os

struct MakerCPP
{
pub mut:
	cxx string
}


fn (mut this MakerCPP) process(states States)
{
	this.cxx = os.getenv_opt("CXX") or { "g++" }
	this.cxx = os.find_abs_path_of_executable(this.cxx) or { os.abs_path(this.cxx) }
	mut process := os.new_process(this.cxx)
	oflags := parse_oflags(states.cflags)
	mut args := ["-o", states.out_path, "-x", "c++", "-c", "-"]
	args << oflags

	process.set_args(args)
	process.set_redirect_stdio()
	println("MakeCPP : starting ${this.cxx}")
	process.run()
	println("MakeCPP : ${this.cxx} startup success ( PID ${process.pid} ), C writing source header...")
	
	process.stdin_write("/** Generated by objbinpack - no one gonna read it this though since this is directly pushed to compiler via stdin */\r")
	process.stdin_write("#include <cstdint>\r\n\n")

	for input in states.inputs {
		varname := input.variable_name 
		process.stdin_write("namespace ${varname} {\n")
		process.stdin_write("\t[[gnu::used]] extern const uint8_t data[];\n\t\t");
		process.stdin_write("\t[[gnu::used]] extern const std::size_t length;\n")
		process.stdin_write("};\n\n")
	}

	for input in states.inputs {
		println("MakeCPP : writing \"${input.file_path}\" as \"${input.variable_name}\"")
		varname := input.variable_name 
		fsize := os.file_size(input.file_path)
		process.stdin_write("\tconst uint8_t ${varname}::data[] = {\n\t\t");
		
		file := os.open(input.file_path)  or { panic(err) }
		mut bytes_read := 0;
		mut buffer := []u8{len:64}
		for !file.eof() {
			buf_read := file.read(mut buffer) or { panic(err) }
			for i in 0 .. buf_read {
				a_byte := buffer[i]
				process.stdin_write("0x${a_byte.hex()}")
				if bytes_read < fsize - 1 {
					process.stdin_write(",")
				}
				bytes_read++
			}
		}

		process.stdin_write("\n\t};\n")

		process.stdin_write("\tconst std::size_t ${varname}::length = ${fsize};\n")
	}

	println("MakeCPP : finishing up")
	os.fd_close(process.stdio_fd[0])
	s_stdout := process.stdout_slurp()
	s_stderr := process.stderr_slurp()
	println("MakeCPP : waiting for ${this.cxx} to exit...")
	process.wait()
	println("${this.cxx} STDOUT: ")
	println(s_stdout)
	println("${this.cxx} STDERR: ")
	println(s_stderr)
	println("MakeCPP : ${this.cxx} exited with code ${process.code} (${process.err}), cleaning up...")
	process.close()
}